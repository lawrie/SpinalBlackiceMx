// Generator : SpinalHDL v1.3.5    git head : f0505d24810c8661a24530409359554b7cfa271a
// Date      : 06/11/2019, 16:39:57
// Component : BlueLed


module BlueLed (
      output  io_blueLed);
  assign io_blueLed = (! 1'b1);
endmodule

